module top_module (
    input clk,
    input reset,
    input [7:0] d,
    output [7:0] q
);

    always@(negedge clk)
        q <= reset ? 6'h0x34 : d;
endmodule
