module top_module ( 
    input clk, 
    input [7:0] d, 
    input [1:0] sel, 
    output [7:0] q 
);

    wire [7:0] q1,q2,q3;
    my_dff8 dflop  (clk,d, q1); 
    my_dff8 dflop1 (clk,q1,q2); 
    my_dff8 dflop2 (clk,q2,q3); 
    
    always@(q3,q1,q2,d,sel) begin  // This is a combinational circuit
     case(sel) 
         4'b0000 : q = d;
         4'b0001 : q = q1;
         4'b0010 : q = q2;
         4'b0011 : q = q3;
     endcase
    end 
endmodule
